`define BLOCK_INSTR_FORMAT_A 0
`define BLOCK_INSTR_FORMAT_B 1

`define BLOCK_INSTR_NOP 			0
`define BLOCK_INSTR_ADD 			1
`define BLOCK_INSTR_SUB 			2
`define BLOCK_INSTR_LSH 			3
`define BLOCK_INSTR_RSH 			4
`define BLOCK_INSTR_ARSH 			5
`define BLOCK_INSTR_MUL 			6
`define BLOCK_INSTR_MADD			7
`define BLOCK_INSTR_ABS				8
`define BLOCK_INSTR_LUT				9
`define BLOCK_INSTR_DELAY_READ 		11
`define BLOCK_INSTR_DELAY_WRITE 	12
`define BLOCK_INSTR_SAVE 			13
`define BLOCK_INSTR_LOAD			14
`define BLOCK_INSTR_MOV				15
`define BLOCK_INSTR_CLAMP			16
`define BLOCK_INSTR_MACZ			17
`define BLOCK_INSTR_MAC				18
`define BLOCK_INSTR_MOV_ACC			19
`define BLOCK_INSTR_LINTERP			20
`define BLOCK_INSTR_FRAC_DELAY		21
`define BLOCK_INSTR_LOAD_ACC		22
`define BLOCK_INSTR_SAVE_ACC		23
`define BLOCK_INSTR_ACC				24
`define BLOCK_INSTR_CLEAR_ACC		25
`define BLOCK_INSTR_MOV_UACC		26

`define BLOCK_OP_TYPE_WIDTH 3

`define BLOCK_INSTR_WIDTH 		32

`define BLOCK_INSTR_OP_WIDTH 	5
`define BLOCK_REG_ADDR_WIDTH   	4
`define BLOCK_PMS_WIDTH			5
`define BLOCK_RES_ADDR_WIDTH	8

`define SHIFT_WIDTH   `BLOCK_PMS_WIDTH

`define N_INSTR_BRANCHES 	4

`define INSTR_BRANCH_MAIN   0
`define INSTR_BRANCH_DELAY  1
`define INSTR_BRANCH_LUT 	2
`define INSTR_BRANCH_MEM 	3
