`define ENGINE_STATE_READY 				0
`define ENGINE_STATE_PROCESSING_WAIT 	1
`define ENGINE_STATE_PROCESSING 		2
`define ENGINE_STATE_MIXING				3