`define CORE_STATE_READY 				0
`define CORE_STATE_BLOCK_START			1
`define CORE_STATE_FETCH_SRC_A			2
`define CORE_STATE_FETCH_SRC_A_2		3
`define CORE_STATE_FETCH_SRC_B			5
`define CORE_STATE_FETCH_SRC_B_2		6
`define CORE_STATE_FETCH_SRC_C			7
`define CORE_STATE_FETCH_SRC_C_2		8
`define CORE_STATE_FINISH_BLOCK			10
`define CORE_STATE_CONTINUE				11
`define CORE_STATE_DISPATCH				12
`define CORE_STATE_FINISH				13
`define CORE_STATE_COMMAND				14

`define CORE_STATE_ADD_1 		110
`define CORE_STATE_ADD_2 		210
`define CORE_STATE_SUB_1 		120
`define CORE_STATE_SUB_2 		220
`define CORE_STATE_MUL_1 		160
`define CORE_STATE_MUL_2 		260
`define CORE_STATE_MAC_1		170
`define CORE_STATE_MAC_2		270
`define CORE_STATE_MAC_3		370
`define CORE_STATE_MAC_4		470
`define CORE_STATE_LUT_1		1100
`define CORE_STATE_ENVD_1 		1110
`define CORE_STATE_DELAY_1 		1120
`define CORE_STATE_GW_1 		1130
`define CORE_STATE_GW_2 		2130
`define CORE_STATE_MOV_1 		1140
`define CORE_STATE_CLAMP_1 		1150
