`define BLOCK_INSTR_NOP 	0
`define BLOCK_INSTR_ADD 	1
`define BLOCK_INSTR_SUB 	2
`define BLOCK_INSTR_LSH 	3
`define BLOCK_INSTR_RSH 	4
`define BLOCK_INSTR_ARSH 	5
`define BLOCK_INSTR_MUL 	6
`define BLOCK_INSTR_MAC		7
`define BLOCK_INSTR_ABS		8
`define BLOCK_INSTR_BIQ_DF1	9
`define BLOCK_INSTR_LUT		10
`define BLOCK_INSTR_ENVD 	11
`define BLOCK_INSTR_DELAY 	12

`define BLOCK_OP_TYPE_WIDTH 3

// Note: ensure 4 * `BLOCK_REG_ADDR_WIDTH + `BLOCK_INSTR_OP_WIDTH + 3 < `BLOCK_INSTR_WIDTH
// and max($clog2(n_channels), $clog2(n_registers)) <= `BLOCK_REG_ADDR_WIDTH
`define BLOCK_INSTR_WIDTH 		32

`define BLOCK_INSTR_OP_WIDTH 	5
`define BLOCK_REG_ADDR_WIDTH   	4
`define BLOCK_PMS_WIDTH			5

// Block FSM states

`define BLOCK_STATE_BEGIN 		0
`define BLOCK_STATE_DONE		1

`define BLOCK_STATE_ADD_WAIT	2
`define BLOCK_STATE_ADD_STORE	3

`define BLOCK_STATE_SUB_WAIT	2
`define BLOCK_STATE_SUB_STORE	3

`define BLOCK_STATE_MUL_WAIT	2
`define BLOCK_STATE_MUL_STORE	3

`define BLOCK_STATE_MAC_MUL_WAIT	2
`define BLOCK_STATE_MAC_ADD_WAIT	3
`define BLOCK_STATE_MAC_STORE		4

`define BLOCK_STATE_BIQUAD_DF1_MUL_1_WAIT 		1

`define BLOCK_STATE_BIQUAD_DF1_MAC_1_MUL_WAIT 	2
`define BLOCK_STATE_BIQUAD_DF1_MAC_1_ACCUMULATE 	3
`define BLOCK_STATE_BIQUAD_DF1_MAC_1_STORE 		4

`define BLOCK_STATE_BIQUAD_DF1_MAC_2_MUL_WAIT 	5
`define BLOCK_STATE_BIQUAD_DF1_MAC_2_ACCUMULATE 	6
`define BLOCK_STATE_BIQUAD_DF1_MAC_2_STORE 		7

`define BLOCK_STATE_BIQUAD_DF1_MAC_3_MUL_WAIT 	8
`define BLOCK_STATE_BIQUAD_DF1_MAC_3_ACCUMULATE 	9
`define BLOCK_STATE_BIQUAD_DF1_MAC_3_STORE 		10

`define BLOCK_STATE_BIQUAD_DF1_MAC_4_MUL_WAIT 	11
`define BLOCK_STATE_BIQUAD_DF1_MAC_4_ACCUMULATE	12
`define BLOCK_STATE_BIQUAD_DF1_SATURATE 		13
`define BLOCK_STATE_BIQUAD_DF1_STORE 			14

`define BLOCK_STATE_LUT_WAIT1 1
`define BLOCK_STATE_LUT_WAIT2 2

`define BLOCK_STATE_ENVD_MUL_1_WAIT 1
`define BLOCK_STATE_ENVD_MUL_2_WAIT 2
`define BLOCK_STATE_ENVD_ADD_WAIT	3
`define BLOCK_STATE_ENVD_STORE		4

`define BLOCK_STATE_DELAY_READ_WAIT 	1
`define BLOCK_STATE_DELAY_MUL_WAIT		2
`define BLOCK_STATE_DELAY_ADD_WAIT		3
`define BLOCK_STATE_DELAY_WRITE_WAIT	4
