`default_nettype none

module top #(
		parameter n_blocks 			= 255,
		parameter data_width 		= 16,
		parameter spi_fifo_length	= 16
	) (
		`ifndef verilator
		input wire crystal,
		`else
		input wire sys_clk,
		`endif

		input  wire cs,
		input  wire mosi,
		output wire miso,
		input  wire sck,

		output wire led0,
		output wire led1,
		output wire led2,
		output wire led3,
		output wire led4,
		output wire led5,

		output wire mclk_out,
		output wire bclk_out,
		output wire lrclk_out,
		
		input  wire i2s_din,
		output wire i2s_dout,

		output wire codec_en
	);
	
	/**********/
	/* Engine */
	/**********/
	
	dsp_engine #(
		.n_blocks(n_blocks),
		.data_width(data_width),
		.spi_fifo_length(spi_fifo_length)
	) engine (
		.clk(sys_clk),
		.reset(reset),

		.in_sample(sample_in),
		.out_sample(sample_out),
	
		.sample_valid(sample_valid),
	
		.command_in(spi_in),
		.command_in_valid(spi_in_valid),

		.current_pipeline(current_pipeline),
		
		.out(out),
		.spi_byte_out(spi_byte_out)
	);
	
	wire [7:0] out;
	wire [7:0] spi_byte_out;
	
	wire current_pipeline;
	
	wire reset = ~pll_lock;
	
	/***********/
	/*   I/O   */
	/***********/

	// Useful LED indicators (active low)
	assign led0 = ~current_pipeline;
	assign led1 = ~out[0];
	assign led3 = ~out[1];
	assign led4 = ~out[2];
	assign led5 = ~out[3];

	// I2S
	wire sample_valid;

	wire [data_width - 1 : 0] sample_out;
	wire [data_width - 1 : 0] sample_in;

	i2s_trx #(.sample_size(data_width)) i2s_driver (
		.sys_clk(sys_clk), .bclk(bclk), .lrclk(lrclk), .din(i2s_din), .dout(i2s_dout),
		.enable(1'b1), .reset(reset), .rx_valid(sample_valid),
		.tx_l(sample_out), .tx_r(sample_out),
		.rx_l(sample_in), .rx_r()
	);
	
	// SPI
	wire [7:0] spi_in;
	wire spi_in_valid;
	
	reg  [4:0] spi_byte_ctr = 0;

	sync_spi_slave spi (
		.clk(sys_clk),
		.reset(reset),

		.sck(sck),
		.cs(cs),
		.mosi(mosi),
		.miso(miso),
		.miso_byte(spi_byte_out),

		.enable(1),

		.mosi_byte(spi_in),
		.data_valid(spi_in_valid)
	);
	
	// Enable power supply to codec when PLL is locked
	assign codec_en = pll_lock;
	
	/**********/
	/* Clocks */
	/**********/
	
	`ifndef verilator // Non-simulated; use crystal and PLL
	wire sys_clk;
	wire pll_lock;
	
	/* PLL to generate main clock from crystal */
	Gowin_rPLL pll(
		.clkout(sys_clk),
		.clkin(crystal),
		.lock(pll_lock)
	);
	`else // Simulated; clock is generated by simulator
	reg pll_lock = 0;
	
	always @(posedge sys_clk)
		pll_lock <= 1;
	`endif

	/* I2S clocks */
	reg mclk = 1'b0;
	reg bclk = 1'b0;
	wire lrclk;
	
	reg [2:0] mclk_ctr = 0;
	reg [3:0] bclk_counter = 4'd0;
	
	reg [5:0] lrclk_counter = 6'd0;
	assign lrclk = lrclk_counter[5];
	
	assign mclk_out  = mclk;
	assign bclk_out  = bclk;
	assign lrclk_out = lrclk;
	
	always @(posedge sys_clk) begin
		if (pll_lock) begin
			if (mclk_ctr == 4) begin
				mclk <= ~mclk;
				mclk_ctr <= 0;

				bclk_counter <= bclk_counter + 1'b1;
				if (bclk_counter == 1) begin
					bclk <= ~bclk;
					bclk_counter <= 0;

					if (bclk)
						lrclk_counter <= lrclk_counter + 1;
					end
			end else begin
				mclk_ctr <= mclk_ctr + 1;
			end
		end   
	end
endmodule

`default_nettype wire
